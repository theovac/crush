library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity sprite_rom is
port 
(	vCounter : in std_logic_vector(8 downto 0);
	pointer : in std_logic_vector(2 downto 0);
	output : out std_logic_vector(39 downto 0)
);
end sprite_rom;

architecture sprite of sprite_rom is
	signal row : std_logic_vector(8 downto 0);
	signal address : std_logic_vector(8 downto 0);

begin

process (vCounter)
begin
	if unsigned(vCounter) < 40 then
		row <= vCounter;
	elsif unsigned(vCounter) < 80 then
		row <= unsigned(vCounter) - 40;
	elsif unsigned(vCounter) <120 then
		row <= unsigned(vCounter) - 80;
	elsif unsigned(vCounter) <160 then
		row <= unsigned(vCounter) - 120;
	elsif unsigned(vCounter) <200 then
		row <= unsigned(vCounter) -160;
	elsif unsigned(vCounter) <240 then
		row <= unsigned(vCounter) -200;
	elsif unsigned(vCounter) <280 then
		row <= unsigned(vCounter) -240;
	elsif unsigned(vCounter) <320 then
		row <= unsigned(vCounter) -280;
	elsif unsigned(vCounter) <360 then
		row <= unsigned(vCounter) -320;
	elsif unsigned(vCounter) <400 then
		row <= unsigned(vCounter) -360;
	elsif unsigned(vCounter) <440 then
		row <= unsigned(vCounter) -400;
	elsif unsigned(vCounter) <480 then
		row <= unsigned(vCounter) -440;
	else 
		row <= (others => '0');
	end if;
end process;


					


address(8 downto 6) <= pointer;
address(5 downto 0) <= row(5 downto 0);


process(address)
begin
case address is

--first sprite icon

when "000000000" => output <= "1111111111111111111111111111111111111111";
when "000000001" => output <= "1000000000000000000000000000000000000001";
when "000000010" => output <= "1000000000000000000000000000000000000001";
when "000000011" => output <= "1000000000000000000000000000000000000001";
when "000000100" => output <= "1000000000000000000000000000000000000001";
when "000000101" => output <= "1000000000000000000000000000000000000001";
when "000000110" => output <= "1000000000000000000000000000000000000001";
when "000000111" => output <= "1000000000000000000000000000000000000001";
when "000001000" => output <= "1000000000000000000000000000000000000001";
when "000001001" => output <= "1000000000000000000000000000000000000001";
when "000001010" => output <= "1000000000000000000000000000000000000001";
when "000001011" => output <= "1000000000000000000000000000000000000001";
when "000001100" => output <= "1000000000000000000000000000000000000001";
when "000001101" => output <= "1000000000000000000000000000000000000001";
when "000001110" => output <= "1000000000000000000000000000000000000001";
when "000001111" => output <= "1000000000000000000000000000000000000001";
when "000010000" => output <= "1000000000000000000000000000000000000001";
when "000010001" => output <= "1000000000000000000000000000000000000001";
when "000010010" => output <= "1000000000000000000000000000000000000001";
when "000010011" => output <= "1000000000000000000000000000000000000001";
when "000010100" => output <= "1000000000000000000000000000000000000001";
when "000010101" => output <= "1000000000000000000000000000000000000001";
when "000010110" => output <= "1000000000000000000000000000000000000001";
when "000010111" => output <= "1000000000000000000000000000000000000001";
when "000011000" => output <= "1000000000000000000000000000000000000001";
when "000011001" => output <= "1000000000000000000000000000000000000001";
when "000011010" => output <= "1000000000000000000000000000000000000001";
when "000011011" => output <= "1000000000000000000000000000000000000001";
when "000011100" => output <= "1000000000000000000000000000000000000001";
when "000011101" => output <= "1000000000000000000000000000000000000001";
when "000011110" => output <= "1000000000000000000000000000000000000001";
when "000011111" => output <= "1000000000000000000000000000000000000001";
when "000100000" => output <= "1000000000000000000000000000000000000001";
when "000100001" => output <= "1000000000000000000000000000000000000001";
when "000100010" => output <= "1000000000000000000000000000000000000001";
when "000100011" => output <= "1000000000000000000000000000000000000001";
when "000100100" => output <= "1000000000000000000000000000000000000001";
when "000100101" => output <= "1000000000000000000000000000000000000001";
when "000100110" => output <= "1000000000000000000000000000000000000001";
when "000100111" => output <= "1111111111111111111111111111111111111111";

--second sprite icon

when "001000000" => output <= "1111111111111111111111111111111111111111";
when "001000001" => output <= "1000000000000000000000000000000000000001";
when "001000010" => output <= "1000000000000000000000000000000000000001";
when "001000011" => output <= "1000000000000000000000000000000000000001";
when "001000100" => output <= "1000000000000000000000000000000000000001";
when "001000101" => output <= "1000000000000000000000000000000000000001";
when "001000110" => output <= "1000000000000000000000000000000000000001";
when "001000111" => output <= "1000000000000000000000000000000000000001";
when "001001000" => output <= "1000000011111111111111111111111100000001";
when "001001001" => output <= "1000000011111111111111111111111100000001";
when "001001010" => output <= "1000000011111111111111111111111100000001";
when "001001011" => output <= "1000000011111111111111111111111100000001";
when "001001100" => output <= "1000000011111111111111111111111100000001";
when "001001101" => output <= "1000000011111111111111111111111100000001";
when "001001110" => output <= "1000000011111111111111111111111100000001";
when "001001111" => output <= "1000000011111111111111111111111100000001";
when "001010000" => output <= "1000000011111111111111111111111100000001";
when "001010001" => output <= "1000000011111111111111111111111100000001";
when "001010010" => output <= "1000000011111111111111111111111100000001";
when "001010011" => output <= "1000000011111111111111111111111100000001";
when "001010100" => output <= "1000000011111111111111111111111100000001";
when "001010101" => output <= "1000000011111111111111111111111100000001";
when "001010110" => output <= "1000000011111111111111111111111100000001";
when "001010111" => output <= "1000000011111111111111111111111100000001";
when "001011000" => output <= "1000000011111111111111111111111100000001";
when "001011001" => output <= "1000000011111111111111111111111100000001";
when "001011010" => output <= "1000000011111111111111111111111100000001";
when "001011011" => output <= "1000000011111111111111111111111100000001";
when "001011100" => output <= "1000000011111111111111111111111100000001";
when "001011101" => output <= "1000000011111111111111111111111100000001";
when "001011110" => output <= "1000000011111111111111111111111100000001";
when "001011111" => output <= "1000000011111111111111111111111100000001";
when "001100000" => output <= "1000000000000000000000000000000000000001";
when "001100001" => output <= "1000000000000000000000000000000000000001";
when "001100010" => output <= "1000000000000000000000000000000000000001";
when "001100011" => output <= "1000000000000000000000000000000000000001";
when "001100100" => output <= "1000000000000000000000000000000000000001";
when "001100101" => output <= "1000000000000000000000000000000000000001";
when "001100110" => output <= "1000000000000000000000000000000000000001";
when "001100111" => output <= "1111111111111111111111111111111111111111";


-- third sprite icon

when "010000000" => output <= "1111111111111111111111111111111111111111";
when "010000001" => output <= "1000000000000000000000000000000000000001";
when "010000010" => output <= "1000000000000000000000000000000000000001";
when "010000011" => output <= "1000000000000000000000000000000000000001";
when "010000100" => output <= "1000000000000000000000000000000000000001";
when "010000101" => output <= "1000000000000000000000000000000000000001";
when "010000110" => output <= "1000000000000000000000000000000000000001";
when "010000111" => output <= "1000000000000000000000000000000000000001";
when "010001000" => output <= "1000000000000011111111111100000000000001";
when "010001001" => output <= "1000000000000011111111111100000000000001";
when "010001010" => output <= "1000000000000011111111111100000000000001";
when "010001011" => output <= "1000000000000011111111111100000000000001";
when "010001100" => output <= "1000000000000011111111111100000000000001";
when "010001101" => output <= "1000000000000011111111111100000000000001";
when "010001110" => output <= "1000000000000011111111111100000000000001";
when "010001111" => output <= "1000000000000011111111111100000000000001";
when "010010000" => output <= "1001111111111111111111111111111111111001";
when "010010001" => output <= "1001111111111111111111111111111111111001";
when "010010010" => output <= "1001111111111111111111111111111111111001";
when "010010011" => output <= "1001111111111111111111111111111111111001";
when "010010100" => output <= "1001111111111111111111111111111111111001";
when "010010101" => output <= "1001111111111111111111111111111111111001";
when "010010110" => output <= "1001111111111111111111111111111111111001";
when "010010111" => output <= "1000000000000011111111111100000000000001";
when "010011000" => output <= "1000000000000011111111111100000000000001";
when "010011001" => output <= "1000000000000011111111111100000000000001";
when "010011010" => output <= "1000000000000011111111111100000000000001";
when "010011011" => output <= "1000000000000011111111111100000000000001";
when "010011100" => output <= "1000000000000011111111111100000000000001";
when "010011101" => output <= "1000000000000011111111111100000000000001";
when "010011110" => output <= "1000000000000011111111111100000000000001";
when "010011111" => output <= "1000000000000011111111111100000000000001";
when "010100000" => output <= "1000000000000000000000000000000000000001";
when "010100001" => output <= "1000000000000000000000000000000000000001";
when "010100010" => output <= "1000000000000000000000000000000000000001";
when "010100011" => output <= "1000000000000000000000000000000000000001";
when "010100100" => output <= "1000000000000000000000000000000000000001";
when "010100101" => output <= "1000000000000000000000000000000000000001";
when "010100110" => output <= "1000000000000000000000000000000000000001";
when "010100111" => output <= "1111111111111111111111111111111111111111";

-- forth sprite icon


when "011000000" => output <= "1111111111111111111111111111111111111111";
when "011000001" => output <= "1000000000000000000000000000000000000001";
when "011000010" => output <= "1000000000000000000000000000000000000001";
when "011000011" => output <= "1000000000000000000000000000000000000001";
when "011000100" => output <= "1000000000000000000000000000000000000001";
when "011000101" => output <= "1000000000000000000000000000000000000001";
when "011000110" => output <= "1000000000000000000000000000000000000001";
when "011000111" => output <= "1000000000000000000000000000000000000001";
when "011001000" => output <= "1000000000000000000110000000000000000001";
when "011001001" => output <= "1000000000000000001111000000000000000001";
when "011001010" => output <= "1000000000000000011111100000000000000001";
when "011001011" => output <= "1000000000000000111111110000000000000001";
when "011001100" => output <= "1000000000000001111111111000000000000001";
when "011001101" => output <= "1000000000000011111111111100000000000001";
when "011001110" => output <= "1000000000000111111111111110000000000001";
when "011001111" => output <= "1000000000001111111111111111000000000001";
when "011010000" => output <= "1000000000011111111111111111100000000001";
when "011010001" => output <= "1000000000111111111111111111110000000001";
when "011010010" => output <= "1000000001111111111111111111111000000001";
when "011010011" => output <= "1000000011111111111111111111111100000001";
when "011010100" => output <= "1000000011111111111111111111111100000001";
when "011010101" => output <= "1000000001111111111111111111111000000001";
when "011010110" => output <= "1000000000111111111111111111110000000001";
when "011010111" => output <= "1000000000011111111111111111100000000001";
when "011011000" => output <= "1000000000001111111111111111000000000001";
when "011011001" => output <= "1000000000000111111111111110000000000001";
when "011011010" => output <= "1000000000000011111111111100000000000001";
when "011011011" => output <= "1000000000000001111111111000000000000001";
when "011011100" => output <= "1000000000000000111111110000000000000001";
when "011011101" => output <= "1000000000000000011111100000000000000001";
when "011011110" => output <= "1000000000000000001111000000000000000001";
when "011011111" => output <= "1000000000000000000110000000000000000001";
when "011100000" => output <= "1000000000000000000000000000000000000001";
when "011100001" => output <= "1000000000000000000000000000000000000001";
when "011100010" => output <= "1000000000000000000000000000000000000001";
when "011100011" => output <= "1000000000000000000000000000000000000001";
when "011100100" => output <= "1000000000000000000000000000000000000001";
when "011100101" => output <= "1000000000000000000000000000000000000001";
when "011100110" => output <= "1000000000000000000000000000000000000001";
when "011100111" => output <= "1111111111111111111111111111111111111111";

--fifth icon

when "100000000" => output <= "1111111111111111111111111111111111111111";
when "100000001" => output <= "1000000000000000000000000000000000000001";
when "100000010" => output <= "1000000000000000000000000000000000000001";
when "100000011" => output <= "1000000000000000000000000000000000000001";
when "100000100" => output <= "1000000000000000000000000000000000000001";
when "100000101" => output <= "1000000000000000000000000000000000000001";
when "100000110" => output <= "1000000000000000000000000000000000000001";
when "100000111" => output <= "1000000000000000000000000000000000000001";
when "100001000" => output <= "1000000000000000000000000000000000000001";
when "100001001" => output <= "1000000000000000000000000000000000000001";
when "100001010" => output <= "1000000000000000000000000000000000000001";
when "100001011" => output <= "1000000000000000000000000000000000000001";
when "100001100" => output <= "1000000000000000000000000000000000000001";
when "100001101" => output <= "1000000000000000000000000000000000000001";
when "100001110" => output <= "1000000000000000000000000000000000000001";
when "100001111" => output <= "1000000000000000000110000000000000000001";
when "100010000" => output <= "1000000000000000001111000000000000000001";
when "100010001" => output <= "1000000000000000011111100000000000000001";
when "100010010" => output <= "1000000000000000111111110000000000000001";
when "100010011" => output <= "1000000000000001111111111000000000000001";
when "100010100" => output <= "1000000000000011111111111100000000000001";
when "100010101" => output <= "1000000000000111111111111110000000000001";
when "100010110" => output <= "1000000000001111111111111111000000000001";
when "100010111" => output <= "1000000000011111111111111111100000000001";
when "100011000" => output <= "1000000000111111111111111111110000000001";
when "100011001" => output <= "1000000001111111111111111111111000000001";
when "100011010" => output <= "1000000011111111111111111111111100000001";
when "100011011" => output <= "1000000111111111111111111111111110000001";
when "100011100" => output <= "1000001111111111111111111111111111000001";
when "100011101" => output <= "1000011111111111111111111111111111100001";
when "100011110" => output <= "1000111111111111111111111111111111110001";
when "100011111" => output <= "1001111111111111111111111111111111111001";
when "100100000" => output <= "1000000000000000000000000000000000000001";
when "100100001" => output <= "1000000000000000000000000000000000000001";
when "100100010" => output <= "1000000000000000000000000000000000000001";
when "100100011" => output <= "1000000000000000000000000000000000000001";
when "100100100" => output <= "1000000000000000000000000000000000000001";
when "100100101" => output <= "1000000000000000000000000000000000000001";
when "100100110" => output <= "1000000000000000000000000000000000000001";
when "100100111" => output <= "1111111111111111111111111111111111111111";

when "101000000" => output <= "1111111111111111111111111111111111111111";
when "101000001" => output <= "1000000000000000000000000000000000000001";
when "101000010" => output <= "1000000000000000000000000000000000000001";
when "101000011" => output <= "1000000000000000000000000000000000000001";
when "101000100" => output <= "1000000000000000000000000000000000000001";
when "101000101" => output <= "1000000000000000000000000000000000000001";
when "101000110" => output <= "1000000000000000000000000000000000000001";
when "101000111" => output <= "1000000000000000000000000000000000000001";
when "101001000" => output <= "1000000000000000000000000000000000000001";
when "101001001" => output <= "1000000000000000000000000000000000000001";
when "101001010" => output <= "1000000111111110000000000000111111000001";
when "101001011" => output <= "1000011111111111100000000111111111110001";
when "101001100" => output <= "1000111111111111110000001111111111111001";
when "101001101" => output <= "1001111111111111111000011111111111111001";
when "101001110" => output <= "1001111111111111111000011111111111111001";
when "101001111" => output <= "1001111111111111111100111111111111111001";
when "101010000" => output <= "1000111111111111111111111111111111110001";
when "101010001" => output <= "1000011111111111111111111111111111100001";
when "101010010" => output <= "1000001111111111111111111111111111000001";
when "101010011" => output <= "1000000111111111111111111111111110000001";
when "101010100" => output <= "1000000011111111111111111111111100000001";
when "101010101" => output <= "1000000001111111111111111111111000000001";
when "101010110" => output <= "1000000000111111111111111111110000000001";
when "101010111" => output <= "1000000000011111111111111111100000000001";
when "101011000" => output <= "1000000000001111111111111111000000000001";
when "101011001" => output <= "1000000000000111111111111110000000000001";
when "101011010" => output <= "1000000000000011111111111100000000000001";
when "101011011" => output <= "1000000000000001111111111000000000000001";
when "101011100" => output <= "1000000000000000111111110000000000000001";
when "101011101" => output <= "1000000000000000011111100000000000000001";
when "101011110" => output <= "1000000000000000001111000000000000000001";
when "101011111" => output <= "1000000000000000000110000000000000000001";
when "101100000" => output <= "1000000000000000000000000000000000000001";
when "101100001" => output <= "1000000000000000000000000000000000000001";
when "101100010" => output <= "1000000000000000000000000000000000000001";
when "101100011" => output <= "1000000000000000000000000000000000000001";
when "101100100" => output <= "1000000000000000000000000000000000000001";
when "101100101" => output <= "1000000000000000000000000000000000000001";
when "101100110" => output <= "1000000000000000000000000000000000000001";
when "101100111" => output <= "1111111111111111111111111111111111111111";

when "110000000" => output <= "1111111111111111111111111111111111111111";
when "110000001" => output <= "1000000000000000000000000000000000000001";
when "110000010" => output <= "1000000000000000000000000000000000000001";
when "110000011" => output <= "1000000000000000000000000000000000000001";
when "110000100" => output <= "1000000000000000000000000000000000000001";
when "110000101" => output <= "1000000000000000000000000000000000000001";
when "110000110" => output <= "1000000000000000000000000000000000000001";
when "110000111" => output <= "1000000000000000000000000000000000000001";
when "110001000" => output <= "1000000000000000011111100000000000000001";
when "110001001" => output <= "1000000000000011111111111100000000000001";
when "110001010" => output <= "1000000000000111111111111110000000000001";
when "110001011" => output <= "1000000000001111111111111111000000000001";
when "110001100" => output <= "1000000000011111111111111111100000000001";
when "110001101" => output <= "1000000000111111111111111111110000000001";
when "110001110" => output <= "1000000001111111111111111111111000000001";
when "110001111" => output <= "1000000001111111111111111111111000000001";
when "110010000" => output <= "1000000001111111111111111111111000000001";
when "110010001" => output <= "1000000011111111111111111111111100000001";
when "110010010" => output <= "1000000011111111111111111111111100000001";
when "110010011" => output <= "1000000011111111111111111111111100000001";
when "110010100" => output <= "1000000011111111111111111111111100000001"; 
when "110010101" => output <= "1000000011111111111111111111111100000001";
when "110010110" => output <= "1000000001111111111111111111111000000001";
when "110010111" => output <= "1000000001111111111111111111111000000001";
when "110011000" => output <= "1000000001111111111111111111111000000001";
when "110011001" => output <= "1000000000111111111111111111110000000001";
when "110011010" => output <= "1000000000011111111111111111100000000001";
when "110011011" => output <= "1000000000001111111111111111000000000001";
when "110011100" => output <= "1000000000000111111111111110000000000001";
when "110011101" => output <= "1000000000000011111111111100000000000001";
when "110011110" => output <= "1000000000000000011111100000000000000001";
when "110011111" => output <= "1000000000000000000000000000000000000001";
when "110100000" => output <= "1000000000000000000000000000000000000001";
when "110100001" => output <= "1000000000000000000000000000000000000001";
when "110100010" => output <= "1000000000000000000000000000000000000001";
when "110100011" => output <= "1000000000000000000000000000000000000001";
when "110100100" => output <= "1000000000000000000000000000000000000001";
when "110100101" => output <= "1000000000000000000000000000000000000001";
when "110100110" => output <= "1000000000000000000000000000000000000001";
when "110100111" => output <= "1111111111111111111111111111111111111111";

when "111000000" => output <= "1111111111111111111111111111111111111111";
when "111000001" => output <= "1000000000000000000000000000000000000001";
when "111000010" => output <= "1000000000000000000000000000000000000001";
when "111000011" => output <= "1000000000000000000000000000000000000001";
when "111000100" => output <= "1000000000000000000000000000000000000001";
when "111000101" => output <= "1000000000000000000000000000000000000001";
when "111000110" => output <= "1000000000000000000000000000000000000001";
when "111000111" => output <= "1000000000000000000000000000000000000001";
when "111001000" => output <= "1000000000000000000000000000000000000001";
when "111001001" => output <= "1000000000000000000000000000000000000001";
when "111001010" => output <= "1000000000000000000000000000000000000001";
when "111001011" => output <= "1000000000000000000000000000000000000001";
when "111001100" => output <= "1000011111111000000000000001111111100001";
when "111001101" => output <= "1000001111111100000000000011111111000001";
when "111001110" => output <= "1000000111111110000000000111111110000001";
when "111001111" => output <= "1000000011111111000000001111111100000001";
when "111010000" => output <= "1000000001111111100000011111111000000001";
when "111010001" => output <= "1000000000111111110000111111110000000001";
when "111010010" => output <= "1000000000011111111001111111100000000001";
when "111010011" => output <= "1000000000001111111111111111000000000001";
when "111010100" => output <= "1000000000000111111111111110000000000001"; --  
when "111010101" => output <= "1000000000001111111111111111000000000001";
when "111010110" => output <= "1000000000011111111001111111100000000001";
when "111010111" => output <= "1000000000111111110000111111110000000001";
when "111011000" => output <= "1000000001111111100000011111111000000001";
when "111011001" => output <= "1000000011111111000000001111111100000001";
when "111011010" => output <= "1000000111111110000000000111111110000001";
when "111011011" => output <= "1000001111111100000000000011111111000001";
when "111011100" => output <= "1000011111111000000000000001111111100001";
when "111011101" => output <= "1000000000000000000000000000000000000001";
when "111011110" => output <= "1000000000000000000000000000000000000001";
when "111011111" => output <= "1000000000000000000000000000000000000001";
when "111100000" => output <= "1000000000000000000000000000000000000001";
when "111100001" => output <= "1000000000000000000000000000000000000001";
when "111100010" => output <= "1000000000000000000000000000000000000001";
when "111100011" => output <= "1000000000000000000000000000000000000001";
when "111100100" => output <= "1000000000000000000000000000000000000001";
when "111100101" => output <= "1000000000000000000000000000000000000001";
when "111100110" => output <= "1000000000000000000000000000000000000001";
when "111100111" => output <= "1111111111111111111111111111111111111111";

when others => output <= "0000000000000000000000000000000000000000";
end case;
end process;
end sprite;

 